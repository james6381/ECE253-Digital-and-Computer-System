module adder(C_in, A, B, C_out, S);
	input C_in;
	input [3:0]A, B;
	output C_out;
	output [3:0]S;
	wire [3:1]C;
	
	full_adder A0(A[0], B[0], C_in, S[0], C[1]);
	full_adder A1(A[1], B[1], C[1], S[1], C[2]);
	full_adder A2(A[2], B[2], C[2], S[2], C[3]);
	full_adder A3(A[3], B[3], C[3], S[3], C_out);
	
endmodule
